module ps2keyb(

	input	wire	clock_50,  	/* 50 мегагерц */
	inout 	wire 	ps2_clock,  /* CLK */
	inout 	wire 	ps2_data,   /* DATA */

);

endmodule
