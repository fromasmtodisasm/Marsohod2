module cpu(

    input  wire        CLK,     // 1.71 МГц
    input  wire        CE,      // Готовность
    output wire [15:0] ADDR,    // Адрес программы или данных
    input  wire [7:0]  DIN,     // Входящие данные
    output reg  [7:0]  DOUT,    // Исходящие данные
    output wire [15:0] EAWR,    // Эффективный адрес для записи
    output reg         WREQ,    // =1 Запись в память по адресу EA
    output reg         RD       // На нисходящем CLK при RD=1, защелка PPU 

);

assign ADDR = AS ? {8'h01, S} : (AM ? EA : PC);
assign EAWR = AS ? {8'h01, S} : EA;

// ---------------------------------------------------------------------

/* Ссылки на микрокод */
`define NDX     5'h01
`define NDY     5'h04
`define ZP      5'h07
`define ZPX     5'h08
`define ZPY     5'h09
`define ABS     5'h0A
`define ABX     5'h0C
`define ABY     5'h0E

// Везде переход к исполнению
`define LAT1    5'h10
`define IMM     5'h11
`define IMP     5'h11
`define ACC     5'h11
`define EXEC    5'h11
`define EXEC2   5'h12
`define EXEC3   5'h13
`define EXEC4   5'h14
// Переход
`define REL     5'h15
`define REL1    5'h16
`define REL2    5'h17
`define LATX    5'h18

initial begin EA = 16'h0000; WREQ = 1'b0; DOUT = 8'h00; RD = 1'b0; end

/* Регистры */
reg  [7:0] A  = 8'h43;
reg  [7:0] X  = 8'h82;
reg  [7:0] Y  = 8'h80;
reg  [7:0] S  = 8'hFF;
reg  [7:0] P  = 8'b00000001;
reg [15:0] PC = 16'h8000;

/* Состояние процессора */
reg         AS     = 1'b0;  /* Указатель стека (приориетнее) */
reg         AM     = 1'b0;  /* 0=PC, 1=EA */
reg  [4:0]  MS     = 3'h0;  /* Исполняемый цикл */
reg  [7:0]  TR     = 3'h0;  /* Temporary Register */
reg  [15:0] EA     = 16'h0000;  /* Эффективный адрес */
reg         WR     = 1'b0;  /* Записать в регистр RA из АЛУ */
reg         FW     = 1'b0;  /* Записать в регистр P из АЛУ */
reg         SW     = 1'b0;  /* Записать в S из АЛУ */
reg         BR     = 1'b0;  /* Если =1, условие выполняется */
reg         ACC    = 1'b0;  /* Указать A вместо DIN */
reg         Cout   = 1'b0;  /* Переносы при вычислении адреса */
reg  [7:0]  opcode = 8'h0;  /* Текущий опкод */
reg         HOP    = 1'b0;  /* =1 Операнду требуется PC++ */
reg  [7:0]  PCL    = 8'h00; /* Для JSR */

/* Некоторые часто употребляемые выражения */
wire [15:0] PCINC   = PC + 1'b1;         /* Инкремент PC */
wire [15:0] PCRel   = PCINC + {{8{DIN[7]}}, DIN[7:0]}; /* Для переходов */
wire [4:0]  MSINC   = MS + 1'b1;         /* Инкремент MS */
wire [15:0] EAINC   = EA + 1'b1;         /* Инкремент EA */
wire [8:0]  XDin    = X + DIN;           /* Для преиндексной адресации */
wire [8:0]  YDin    = Y + DIN;           /* Для постиндексной адресации */
wire [7:0]  HIDin   = DIN + Cout;        /* Перенос */
wire [15:0] EADIN   = {DIN,   TR};
wire [15:0] EADIH   = {HIDin, TR};
wire        INCDEC  = ({opcode[7:6], opcode[2:0]} == 5'b11_1_10) || /* INC/DEC */
                      ({opcode[7],   opcode[2:0]} == 4'b0__1_10);   /* Сдвиговые */

wire        Latency = Cout | (opcode[7:5] == 3'b100) | INCDEC; /* STA, Cout, Сдвиговые */
wire [4:0]  LATAD   = Latency ? `LAT1 : `EXEC; /* Код адреса при Latency */

/* Исполнение микрокода */
always @(posedge CLK) begin

    case (MS)

        /* ИНИЦИАЛИЗАЦИЯ */
        4'h0: begin

            casex (DIN)

                8'bxxx_000_x1: begin MS <= `NDX; HOP <= 1'b1; end // Indirect, X
                8'bxxx_010_x1, // Immediate
                8'b1xx_000_x1: begin MS <= `IMM; HOP <= 1'b1; end
                8'bxxx_100_x1: begin MS <= `NDY; HOP <= 1'b1; end // Indirect, Y
                8'bxxx_110_x1: begin MS <= `ABY; HOP <= 1'b1; end // Absolute, Y
                8'bxxx_001_xx: begin MS <= `ZP;  HOP <= 1'b1; end  // ZeroPage
                8'bxxx_011_xx, // Absolute
                8'b001_000_00: begin MS <= `ABS; HOP <= 1'b1; end
                8'b10x_101_1x: begin MS <= `ZPY; HOP <= 1'b1; end // ZeroPage, Y
                8'bxxx_101_xx: begin MS <= `ZPX; HOP <= 1'b1; end // ZeroPage, X
                8'b10x_111_1x: begin MS <= `ABY; HOP <= 1'b1; end // Absolute, Y
                8'bxxx_111_xx: begin MS <= `ABX; HOP <= 1'b1; end // Absolute, X
                8'bxxx_100_00: begin MS <= `REL; HOP <= 1'b1; end // Relative
                8'b0xx_010_10: begin MS <= `ACC; HOP <= 1'b0; end // Accumulator
                default:       begin MS <= `IMP; HOP <= 1'b0; end

            endcase

            PC      <= PCINC; /* PC++ */
            AS      <= 1'b0;  /* Указатель стека */
            RD      <= 1'b0;  /* Для PPU */
            WREQ    <= 1'b0;  /* Отключение записи в память EA */
            opcode  <= DIN;   /* Принять новый опкод */

        end

        /* АДРЕСАЦИЯ */

        /* Indirect, X */
        // -------------------------------------------------------------
        4'h1: begin MS <= MSINC; EA <= XDin[7:0]; AM <= 1'b1; Cout <= XDin[8]; end
        4'h2: begin MS <= MSINC; EA <= EAINC;     TR <= DIN;  end
        4'h3: begin MS <= `LATX; EA <= EADIN;     RD <= 1'b1; end

        /* Indirect, Y */
        // -------------------------------------------------------------
        4'h4: begin MS <= MSINC; EA <= DIN;   AM <= 1'b1; end
        4'h5: begin MS <= MSINC; EA <= EAINC; TR <= YDin[7:0]; Cout <= YDin[8]; end
        4'h6: begin MS <= LATAD; EA <= EADIH; RD <= 1'b1; end

        /* ZP */
        // -------------------------------------------------------------
        4'h7: begin MS <= `EXEC; EA <= DIN;       RD <= 1'b1; AM <= 1'b1; end

        /* ZP,X */
        // -------------------------------------------------------------
        4'h8: begin MS <= `LAT1; EA <= XDin[7:0]; RD <= 1'b1; AM <= 1'b1; end

        /* ZP,Y */
        // -------------------------------------------------------------
        4'h9: begin MS <= `LAT1; EA <= YDin[7:0]; RD <= 1'b1; AM <= 1'b1; end

        /* Absolute */
        // -------------------------------------------------------------
        4'hA: begin MS <= MSINC; TR <= DIN;    PC <= PCINC;  end
        4'hB: 
        
            /* JMP ABS */
            if (opcode == 8'h4C) 
                 begin PC <= EADIN; MS <= 1'b0; end
            else begin AM <= 1'b1;  MS <= `EXEC; EA <= EADIN; RD <= 1'b1; end
            

        /* Absolute,X */
        // -------------------------------------------------------------
        4'hC: begin MS <= MSINC; TR <= XDin[7:0]; PC <= PCINC; Cout <= XDin[8]; end
        4'hD: begin MS <= LATAD; EA <= EADIH;     RD <= 1'b1;  AM <= 1'b1; end

        /* Absolute,Y */
        // -------------------------------------------------------------
        4'hE: begin MS <= MSINC; TR <= YDin[7:0]; PC <= PCINC; Cout <= YDin[8]; end
        4'hF: begin MS <= LATAD; EA <= EADIH;     RD <= 1'b1;  AM <= 1'b1; end

        /* Отложенный такт (для адресации) */
        `LAT1: MS <= `EXEC;
        
        /* Для (I,X) если X превысил границу ZP */
        `LATX: if (Cout) MS <= `LAT1; else MS <= `EXEC;

        /* Исполнение инструкции */
        // -------------------------------------------------------------

        /* Исполнение инструкции */
        `EXEC: begin

            RD  <= 1'b0;
            PCL <= PC[7:0];

            /* Инкремент PC по завершении разбора адреса */
            if (HOP) PC <= PCINC; 

            casex (opcode)

                /* STA/STY/STX для АЛУ */
                8'b100_xxx_01, 
                8'b100_xx1_x0: {AM, MS, WREQ, DOUT} <= {1'b0, 5'h0,  1'b1, AR[7:0]};
                
                /* JMP Indirect */
                8'b011_011_00: {MS, TR, EA} <= {MSINC, DIN, EA};

                /* ROL/ROR/ASR/LSR/DEC/INC <mem> */
                8'b0xx_xx1_10,
                8'b11x_xx1_10: {AM, MS, WREQ, DOUT} <= {1'b0, MSINC, 1'b1, AR[7:0]};
                
                /* JSR: Записываем в стек */
                8'b001_000_00: {AS, MS, WREQ, DOUT} <= {1'b1, MSINC, 1'b1, PC[15:8]};
                
                /* RTS */
                8'b011_000_00: {AS, MS} <= {1'b1, MSINC};
                
                /* PHP */
                8'b000_010_00: {AS, MS, WREQ, DOUT} <= {1'b1, MSINC, 1'b1, P[7:6], 2'b11, P[3:0]};                
                
                /* PHA */
                8'b010_010_00: {AS, MS, WREQ, DOUT} <= {1'b1, MSINC, 1'b1, A};     
                
                /* PLP, PLA */
                8'b0x1_010_00: {AS, MS} <= {1'b1, MSINC};
                
                // По умолчанию, завершение инструкции
                default: {AM, MS} <= 2'b00;

            endcase

        end
        
        /* Для особых инструкции */
        // -------------------------------------------------------------
        
        `EXEC2: casex (opcode)
        
            8'b001_000_00: begin MS <= MSINC; DOUT <= PCL; end /* JSR */
            8'b011_000_00: begin MS <= MSINC; PC[7:0] <= DIN; end /* RTS */
            8'b011_011_00: begin MS <= 1'b0;  AM <= 1'b0; PC <= EADIN; end /* JMP IND */
            8'b0x0_010_00: begin MS <= 1'b0; {AM, AS, WREQ} <= 3'b000; end /* PHP, PHA */
                  default: begin MS <= MSINC; {AM, AS, WREQ} <= 3'b000; end
        
        endcase
                
        `EXEC3: casex (opcode)
        
            8'b001_000_00: begin MS <= 1'b0; PC <= EA; {AS, WREQ, AM} <= 3'b000; end /* JSR */
            8'b011_000_00: begin MS <= MSINC; PC[15:8] <= DIN; end /* RTS */
                  default: begin MS <= 1'b0; end
                  
        endcase
        
        `EXEC4: casex (opcode)
        
            8'b011_000_00: begin MS <= `REL2; /* +1T */ {AS, AM} <= 2'b00; PC <= PCINC; end /* RTS */
            8'b0x1_010_00: begin MS <= MSINC; AS <= 1'b0; end /* PLP, PLA */
            
        endcase
        

        /* Исполнение инструкции B<cc> */
        // -------------------------------------------------------------

        `REL: begin
        
            if (BR) begin PC <= PCRel; MS <= PCRel[15:8] == PC[15:8] ? `REL2 : `REL1; end
            else    begin PC <= PCINC; MS <= 1'b0; end
    
        end

        `REL1: begin MS <= MSINC; end /* +2T если превышение границ */
        `REL2: begin MS <= 1'b0; end  /* +1T если переход */

    endcase

end

/* Подготовка данных на этапах исполнения */
// ---------------------------------------------------------------------

always @* begin

    alu = {1'b0, opcode[7:5]}; /* По умолчанию */
    RA  = 2'b00; /* A */
    RB  = 2'b00; /* DIN */
    WR  = 1'b0;
    FW  = 1'b0;
    SW  = 1'b0;  /* Stack Write */
    ACC = 1'b0;
    BR  = 1'b0; /* Условие выполнения Branch */

    case (opcode[7:6])
                        
        /* S */ 2'b00: BR = (P[7] == opcode[5]);
        /* V */ 2'b01: BR = (P[6] == opcode[5]);
        /* C */ 2'b10: BR = (P[0] == opcode[5]);
        /* Z */ 2'b11: BR = (P[1] == opcode[5]);
                
    endcase
    
    case (MS)
    `EXEC: casex (opcode)

        /* STA, CMP */
        8'b1x0_xxx_01: FW = opcode[6];

        /* ADC, SBC, AND, ORA, EOR, LDA */
        8'bxxx_xxx_01: {WR, FW} = 2'b11;
        
        /* ROL,ROR,ASL,LSR ACC */
        8'b0xx_010_10: {alu, ACC, RB, RA, FW, WR} = {2'b10, opcode[6:5], 1'b1, 6'b00_00_11};

        /* ASL,ROL,LSR,ROR <mem> */
        8'b0xx_xx1_10: {alu, FW} = {2'b10, opcode[6:5], 1'b1};
        
        /* DEC/INC */
        8'b11x_xx1_10: {alu, FW} = {3'b111, opcode[5], 1'b1};

        /* STY, STX */
        8'b100_xx1_00: {RA} = 2'b10; // Y
        8'b100_xx1_10: {RA} = 2'b01; // X
        
        /* LDY */
        8'b101_xx1_00,
        8'b101_000_00: {WR, RA, FW} = 4'b1_10_1;
        
        /* LDX */
        8'b101_xx1_10,
        8'b101_000_10: {WR, RA, FW} = 4'b1_01_1;
        
        /* CPY */
        8'b110_xx1_00,
        8'b110_000_00: {RA, FW} = 3'b10_1;
        
        /* CPX */
        8'b111_xx1_00,
        8'b111_000_00: {alu, RA, FW} = 7'b0110_01_1;

        /* CLC, SEC, CLI, SEI, CLV, CLD, SED */
        8'bxxx_110_00: {alu, FW} = 5'b1100_1;
        
        /* BIT */
        8'b001_0x1_00: {alu, FW} = 5'b1101_1;
        
        /* Transfer */
        8'b100_010_00: {alu, RA, RB, WR, FW} = 10'b1110_10_10_11; /* DEY */
        8'b110_010_10: {alu, RA, RB, WR, FW} = 10'b1110_01_01_11; /* DEX */
        8'b110_010_00: {alu, RA, RB, WR, FW} = 10'b1111_10_10_11; /* INY */
        8'b111_010_00: {alu, RA, RB, WR, FW} = 10'b1111_01_01_11; /* INX */
                        
        /* TAX, TAY */
        8'b101_010_10: {alu, RB, RA, FW, WR, ACC} = 11'b0101_00_01_111;
        8'b101_010_00: {alu, RB, RA, FW, WR, ACC} = 11'b0101_00_10_111;        
        8'b100_110_10: {alu, RB, SW}     = 8'b0101_01_1;  /* TXS */
        8'b100_110_00: {alu, RB, FW, WR} = 8'b0101_10_11; /* TYA */        
        8'b100_010_10: {alu, RB, FW, WR} = 8'b0101_01_11; /* TXA */        
        8'b101_110_10: {alu, RB, RA, FW, WR} = 10'b0101_11_01_11; /* TSX */
        
        /* RTS, PLP, PLA */
        8'b011_000_00,
        8'b0x1_010_00: {alu, RB, SW} = 7'b1111_11_1; 
        
    endcase
    
    /* Специальные инструкции управления */
    `EXEC2: casex (opcode)
        
        8'b011_000_00: {alu, RB, SW} = 7'b1111_11_1; /* RTS */
        8'b001_000_00,
        8'b0x0_010_00: {alu, RB, SW} = 7'b1110_11_1; /* JSR, PHP, PHA */             
        8'b001_010_00: {RA, WR} = 3'b11_1; /* PLP */
        8'b011_010_00: {RA, WR, alu} = 7'b00_1_0101; /* PLA */
    
    endcase
    
    `EXEC3: casex (opcode)

        /* JSR */
        8'b001_000_00: {alu, RB, SW} = 7'b1110_11_1;
    
    endcase
    
    endcase



end

/* Запись результата */
// ---------------------------------------------------------------------

always @(posedge CLK) begin

    /* Писать результат АЛУ */
    if (WR) case (RA)
        2'b00: A <= AR;
        2'b01: X <= AR;
        2'b10: Y <= AR;
    endcase

    /* Писать флаги */
    if (WR && RA == 2'b11) /* PLP */
        P <= DIN;
    else if (FW)  
        P <= AF;
    
    /* Записать в регистр S результат */
    if (SW) S <= AR;

end

/* Вычислительное устройство */
// ---------------------------------------------------------------------

reg [3:0] alu = 4'h0;
reg [1:0] RA = 2'b00;
reg [1:0] RB = 2'b00;
reg [7:0] Ax;
reg [7:0] Bx;
reg [7:0] AR;
reg [7:0] AF;

always @* begin

    case (RA)
        2'b00: Ax = A;
        2'b01: Ax = X;
        2'b10: Ax = Y;
        2'b11: Ax = 0;
    endcase

    case (RB)
        2'b00: Bx = (ACC ? A : DIN);
        2'b01: Bx = X;
        2'b10: Bx = Y;
        2'b11: Bx = S;
    endcase

end

alu ALU(

    /* Вход */  Ax, Bx, alu, P, opcode[7:5],
    /* Выход */ AR, AF

);

endmodule
