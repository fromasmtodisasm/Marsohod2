module cpu8632();

endmodule
