/*
 * 8-������ ���������
 * 
 * - �� ������ ���������� 6502
 * - �� �������� 25 ���
 */
 
module demo_processor(
   
    // ������������ ���������� �� ����������� ������� 25 ���
    input   wire        clock_25,
    
    // 8-������ ���� ������
    input   wire [7:0]  i_data,         // �������� ������
    output  reg  [15:0] o_addr,         // 16-������ ����� (64 �� �������� ������������)
    output  reg  [7:0]  o_data,         // ������ ��� ������
    output  reg         o_wr            // ������ � ������

);

/*
 * ��������
 */
 
reg [7:0]  a; // �����������
reg [7:0]  x; // ��������� �������
reg [7:0]  y; // ��������� �������
reg [7:0]  p; // �����
reg [7:0]  s; // ���� $100-$1FF
reg [15:0] pc; // ������� ������

/*
 * ���������
 */

reg [3:0] t;    // ������� ��������� ����������

/*
 * ������������� ��������� ��������
 */

initial begin

    a = 8'h00;
    x = 8'h00; y = 8'h00;
    p = 8'h00; s = 8'h00;
    
    t = 4'h0;
    
    // ������ ��������� �������
    pc     = 16'h0000;
    o_addr = 16'h0000;
    
    o_data = 8'h00;
    o_wr = 1'b0;

end

/*
 * ���������� ������
 */
 
// ����������-���������� ���������� [aaaxxx01]
wire c_arithlogic = i_data[1:0] == 2'b01;

/*
 * ������� ������������ ������
 */

always @(posedge clock_25) begin

    case (t)
    
        /*
         * ���������� ������ ���������� ����� ����������
         */
    
        4'h0: begin
        
        end

    endcase

end

endmodule
