module vga(

    // 100 мегагерц
    input   wire        clk,

    // Выходные данные
    output  reg  [4:0]  red,        // 5 бит на красный (4,3,2,1,0)
    output  reg  [5:0]  green,      // 6 бит на зеленый (5,4,3,2,1,0)
    output  reg  [4:0]  blue,       // 5 бит на синий (4,3,2,1,0)
    output  wire        hs,         // синхросигнал горизонтальной развертки
    output  wire        vs,          // синхросигнал вертикальной развертки
    
    output  reg  [11:0] adapter_font,  // 2^12 = 4096 байт
    input   wire [7:0]  adapter_data   // полученные данные от знакогенератора

);

// 640 (видимая область) + 48 (задний порожек) + 96 (синхронизация) + 16 (передний порожек)
// 640 + 48 = [688, 688 + 96 = 784]
assign hs = x >= (640 + 48) && x < 764;

// 480 + 33 + 2 + 10
assign vs = y >= (480 + 33) && y < (480 + 33 + 2);

// В этих регистрах мы будем хранить текущее положение луча на экране
reg [9:0] x = 1'b0; // 2^10 = 1024 точек возможно
reg [9:0] y = 1'b0;

// Объявим регистры со временными данными
reg [7:0] current_char;
reg [7:0] current_data;

// Извлекаем текущий бит (от 0 до 7) в зависимости от положения луча x
wire current_bit = current_data[ x[2:0] ];

// 2х битный счетчик
reg [1:0] clock_divider;

// Делитель частоты. На входе частота - 100 мгц, а на выходе будет 25 Мгц
always @(posedge clk) clock_divider <= clock_divider + 1'b1;

// Когда бит 1 переходит из состояния 0 в состояние 1, это значит, что
// будет осциллироваться на частоте 25 мгц (в 4 раза медленее, чем 100 мгц)
always @(posedge clock_divider[1]) begin

    // аналогично этой конструции на C
    // if (x == 799) x = 0; else x += 1;
    x <= x == 10'd799 ? 1'b0 : (x + 1'b1);
    
    // Когда достигаем конца горизонтальной линии, переходим к Y+1
    if (x == 10'd799) begin
    
        // if (x == 524) y = 0; else y += 1;
        y <= y == 10'd524 ? 1'b0 : (y + 1'b1);

    end
    
    // Мы находимся в видимой области рисования
    if (x < 640 && y < 480) begin
    
        // 640 / 80 = 8
        case (x[2:0])
        
            // пусть пока экран заполнится буквой A
            3'b001: current_char <= 8'h41;  
            
            // Делаем запрос на поиск части символа
            // {current_char, y[3:0]} = current_char * 16 + (y % 16)
            3'b110: adapter_font <= {current_char, y[3:0]};
            
            // Читаем ответ от знакогенератора (через 4 такта на скорости 100 мгц)
            // Или через 1 такт на скорости 25 Мгц, на которой мы сейчас и работаем
            3'b111: current_data <= adapter_data;

        endcase
    
        // Если текущий рисуемый бит =1, то рисовать белым цветом
        // Слегка сероватый фон надо сделать, чтобы меня понял монитор
        red   <= current_bit ? 5'h1F : 5'h03;
        green <= current_bit ? 6'h3F : 6'h03;
        blue  <= current_bit ? 5'h1F : 5'h03;
    
    // В невидимой области мы ДОЛЖНЫ очищать в черный цвет
    // иначе видеоадаптер работать будет неправильно
    end else begin
    
        red   <= 1'b0;
        green <= 1'b0;
        blue  <= 1'b0;
    
    end

end

endmodule
