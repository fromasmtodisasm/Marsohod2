/* 
 * Не находится в ведении копирайтов. Сделан, как кофе с утра.
 * Реклама: я кот, хозяин спит, лей вискаса, а то разодру обои.
 */
 
module z80(

    // О`клок
    input wire          clk,    /* 25 Мгц. Любой. */

    // Кот    #1 Порт
    output reg [15:0]   Ca,     /* Адрес памяти для считывания кода */
    input wire [7:0]    Ci,     /* Считанный код */
    
    // Данные #2 Порт
    output reg [15:0]   Da,     /* Для считывания данных */
    input wire [7:0]    Di,     /* Считанные данные */
    output reg [7:0]    Do,     /* Данные на запись */
    output reg          Dw      /* Сигнал записи */

);

// ---------------------------------------------------------------------
/* Основной набор регистров (8x8 = 256 бит) */
reg [7:0]  B; reg [7:0] C;
reg [7:0]  D; reg [7:0] E;
reg [7:0]  H; reg [7:0] L;
reg [7:0]  A; reg [7:0] F;
reg [15:0] IX;
reg [15:0] IY;
reg [15:0] SP;
reg [15:0] PC;

/* Дополнительный набор. Регистры много занимают памяти в ПЛИС. */
reg [7:0] B_; reg [7:0] C_;
reg [7:0] D_; reg [7:0] E_;
reg [7:0] H_; reg [7:0] L_;
reg [7:0] A_; reg [7:0] F_;

/* Текущий регистр */
reg [2:0] Rq;   /* Запрос чтения */
reg [7:0] Rc;   /* Ответ чтения */

/* Для записи в регистр */
reg [2:0] Wn;   /* Номер регистра */
reg [7:0] Wo;   /* Значение */
reg       We;   /* Сигнал записи на следующем такте */

/* Префиксирование */
reg [1:0] Px;   /* Префиксировано 00 - HL; 01 - IX; 10 - IY; 11 - ?? */
reg [7:0] Hp;   /* Регистр H */
reg [7:0] Lp;   /* Регистр L */

// Состояние процессора
// ---------------------------------------------------------------------
reg [1:0] M_cycle;

// ---------------------------------------------------------------------

/* Инициализация регистров */
initial begin

    PC   = 16'h0000;
    SP   = 16'h0000;
    IX   = 16'h0000;
    IY   = 16'h0000;
    
    Rq   = 3'b000;
    Px   = 2'b00;
    T    = 8'h00;
    
    M_cycle = 1'b0;
    
    //                                      B      C      D      E      H      L      A      F
    {B,  C,  D,  E,  H,  L,  A,  F } = {8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h25, 8'h00};
    {B_, C_, D_, E_, H_, L_, A_, F_} = {8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFA, 8'h00};

end

// Эмуляция микрокода
// ---------------------------------------------------------------------

reg [1:0]   mPCinc;           /* Увеличить PC + mPCinc на следующем такте */

reg         mPCrel;           /* Если =1, переход на jmpRel */
reg         mPCjmp;           /* Признак, что есть переход на PCtmp */
reg [15:0]  PCrel;            /* Вычисление относительн PC перехода 8 бит */

reg         mCycleInc;        /* Увеличить M_cycle */
reg         mEXAF;            /* На следующем такте развернуть AF, AF' */
reg         mBDec;            /* B = B - 1 */

reg [1:0]   mWe16;            /* Запись в 16-битный регистр Wn[1:0] */
reg [1:0]   mT;               /* Действия с регистром T */
reg [7:0]   T;                /* Временное значение */

/* Кеш опкода между M_cycle */
reg [7:0]   opcache;      

/* Источник опкода */
wire [7:0]  opcode = (M_cycle == 1'b0) ? Ci : opcache;  

/* Проверка условий */
wire [3:0]  condition = { F[7], F[2], F[6], F[0] };

// ---------------------------------------------------------------------

always @* begin

    Ca          = PC;
    Da          = PC + 1'b1; /* Ускорение чтения инструкции */
    Dw          = 1'b0;
    
    /* Секция переходов */
    mPCinc      = 2'b01;
    mPCjmp      = 1'b0;
    mPCrel      = 1'b0;      
     PCrel      = PC + {{8{Di[7]}}, Di[7:0]} + 2'h2;
    
    mCycleInc   = 1'b0;
    mEXAF       = 1'b0;
    mT          = 2'b00;
    Wn          = opcode[5:3];
    mWe16       = 2'b00;

    casex (opcode)
    
        // 1T NOP
        8'b00_000_000: begin /* NOP */ end
        
        // 1T EX AF, AF'
        8'b00_001_000: mEXAF = 1'b1; 
        
        // 1T DJNZ *
        8'b00_010_000: {mBDec, mPCinc, mPCrel} = {1'b1, 2'b10, (B != 8'h00) };

        // 1T JR *
        8'b00_011_000: {mPCrel} = {1'b1};
        
        // 1T JR {NC, C, NZ, Z}, *
        8'b00_1xx_000: {mPCinc, mPCrel} = {2'b10, condition[ opcode[4] ] == opcode[3] };
        
        // 2T LD r16, **
        8'b00_xx0_001: case (M_cycle)
        
            /* Запись из Di -> T[7:0], PC += 2 */
            1'b0: {mCycleInc, mT} = {1'b1, 2'b01};
            
            /* Запись {Di, T[7:0]} -> r16 */
            1'b1: {mWe16, Wn[1:0]} = {2'b01, opcode[5:4]};
        
        endcase
    
    endcase

end

// Тактирование. Основная логика
// ---------------------------------------------------------------------

always @(posedge clk) begin

    /* Переходы */
    PC <= mPCrel ? PCrel :  PC + mPCinc;
    
    /* Запись опкода в кеш */
    if (M_cycle == 1'b0)
        opcache <= Ci;
        
    /* Обработка T16 */
    case (mT)
        2'b01: T[7:0] <= Di;
    endcase    
    
    /* Сброс, если последний опкод, либо финализировать */
    M_cycle <= (mCycleInc ? M_cycle + 1'b1 : 1'b0);

end

// Выборка регистра
// ---------------------------------------------------------------------

/* Чтение из регистров */
always @(Rq, Px, mEXAF) begin

    case (Px)
        2'b00: begin Hp = H;        Lp = L; end
        2'b01: begin Hp = IX[15:8]; Lp = IX[7:0]; end
        2'b10: begin Hp = IY[15:8]; Lp = IY[7:0]; end
    endcase
        
    /* Другие инструкции */
    case (Rq)
        
        3'b000: Rc = B;  3'b001: Rc = C;
        3'b010: Rc = D;  3'b011: Rc = E;
        3'b100: Rc = Hp; 3'b101: Rc = Lp;
        3'b110: Rc = Di; 3'b111: Rc = A; 
    
    endcase

end

/* Запись в регистры */
always @(posedge clk) begin

    /* Команда EX AF, AF' */
    if (mEXAF) {A, A_, F, F_} <= {A_, A, F_, F};
    
    /* Уменьшение B = B - 1 */
    else if (mBDec) B <= B - 1'b1;    
    
    /* Запись в регистр 16 бит из памяти {Di, T[7:0]} */
    else if (mWe16 == 2'b01) begin
    
        case (Wn[1:0])
        
            2'b00: {B, C} <= {Di, T[7:0]};
            2'b01: {D, E} <= {Di, T[7:0]};
            2'b10: {H, L} <= {Di, T[7:0]};
            2'b11: SP     <= {Di, T[7:0]};

        endcase
    
    end
        
    /* Регистр */
    else if (We) begin

        case (Wn)
            3'b000: B <= Wo;  3'b001: C <= Wo;
            3'b010: D <= Wo;  3'b011: E <= Wo;
            3'b100: case (Px) 2'b00:  H <= Wo; 2'b01: IX[15:8] <= Wo; 2'b10: IY[15:8] <= Wo; endcase
            3'b101: case (Px) 2'b00:  L <= Wo; 2'b01: IX[ 7:0] <= Wo; 2'b10: IY[ 7:0] <= Wo; endcase
            // 3'b110: /* Запись в память обрабатывается отдельно */ begin Dw <= We; Do <= Wo;  end
            3'b111: A <= Wo;
        endcase

    end
    
    /* Флаги */
    // ... 
    
    // Другое (SP и прочее)

end

endmodule
