module vga(

    // 100 мегагерц
    input   wire        clk,

    // Выходные данные
    output  reg  [4:0]  red,        // 5 бит на красный (4,3,2,1,0)
    output  reg  [5:0]  green,      // 6 бит на зеленый (5,4,3,2,1,0)
    output  reg  [4:0]  blue,       // 5 бит на синий (4,3,2,1,0)
    output  wire        hs,         // синхросигнал горизонтальной развертки
    output  wire        vs          // синхросигнал вертикальной развертки

);

// 640 (видимая область) + 48 (задний порожек) + 96 (синхронизация) + 16 (передний порожек)
// 640 + 48 = [688, 688 + 96 = 784]
assign hs = x >= (640 + 48) && x < 764;

// 480 + 33 + 2 + 10
assign vs = y >= (480 + 33) && y < (480 + 33 + 2);

// В этих регистрах мы будем хранить текущее положение луча на экране
reg [9:0] x = 1'b0; // 2^10 = 1024 точек возможно
reg [9:0] y = 1'b0;

// 2х битный счетчик
reg [1:0] clock_divider;

// Делитель частоты. На входе частота - 100 мгц, а на выходе будет 25 Мгц
always @(posedge clk) clock_divider <= clock_divider + 1'b1;

// Когда бит 1 переходит из состояния 0 в состояние 1, это значит, что
// будет осциллироваться на частоте 25 мгц (в 4 раза медленее, чем 100 мгц)
always @(posedge clock_divider[1]) begin

    // аналогично этой конструции на C
    // if (x == 799) x = 0; else x += 1;
    x <= x == 10'd799 ? 1'b0 : (x + 1'b1);
    
    // Когда достигаем конца горизонтальной линии, переходим к Y+1
    if (x == 10'd799) begin
    
        // if (x == 524) y = 0; else y += 1;
        y <= y == 10'd524 ? 1'b0 : (y + 1'b1);

    end
    
    // Мы находимся в видимой области рисования
    if (x < 640 && y < 480) begin
    
        // типичная XOR текстура, сейчас заценим...
        red   <= x[4:0] ^ y[4:0]; // 5'h1F;
        green <= x[5:0] ^ y[5:0]; // 6'h3F;
        blue  <= x[4:0] ^ y[4:0]; // 5'h1F;    
    
    // В невидимой области мы ДОЛЖНЫ очищать в черный цвет
    // иначе видеоадаптер работать будет неправильно
    end else begin
    
        red   <= 1'b0;
        green <= 1'b0;
        blue  <= 1'b0;
    
    end

end

endmodule
