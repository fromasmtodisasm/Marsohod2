/*
 * Простой 8-битный процессор
 * 
 * - на основе инструкции 6502
 * - на скорости 25 мгц
 */
 
module processor(
   
    // Тактирование процессора на стандартной частоте 25 Мгц
    input   wire        clock_25,
    
    // 8-битная шина данных
    input   wire [7:0]  i_data,         // Входящие данные
    output  wire [15:0] o_addr,         // 16-битный адрес (64 кб адресное пространство)
    output  reg  [7:0]  o_data,         // Данные для записи
    output  reg         o_wr            // Запись в память

);

/*
 * Роутинг
 */

assign o_addr = alt ? addr : pc;

/*
 * Регистры
 */
 
reg [7:0]  a; // Аккумулятор
reg [7:0]  x; // Индексный регистр
reg [7:0]  y; // Индексный регистр
reg [7:0]  p; // Флаги
reg [7:0]  s; // Стек $100-$1FF
reg [15:0] pc; // Регистр адреса

/*
 * Состояния
 */

reg [3:0]  t;        // Текущее состояние процессора
reg [2:0]  am;       // Address Mode = 0..7, декодирование
reg [7:0]  op_cache; // Предущущее состояние опкода
reg        alt;      // Если =1, то смотрит в память [addr], иначе на [pc]
reg [15:0] addr;     // Указатель на рабочую область памяти
reg [7:0]  tmp8;     // Временный 8-bit регистр

/*
 * Инициализация первичных значений
 */

initial begin

    a = 8'h00;
    x = 8'h00; y = 8'h00;
    p = 8'h00; s = 8'h00;
    
    t = 4'h0;
    am = 3'h0;
    alt = 1'b0;
    
    // Должны совпадать вначале
    pc     = 16'h0000;
    addr   = 16'h0000;
    
    op_cache = 8'h00;
    o_data = 8'h00;
    o_wr = 1'b0;

end

/*
 * Дешифратор кода операции
 */

// Актуальный опкод всё время
wire [7:0] opcode = t ? op_cache : i_data;

/*
 * Главная процессорная логика
 */

always @(posedge clock_25) begin

    case (t)
    
        /* 1. Дешифрация инструкции - выбор режима операнда */   
        4'h0: begin
        
            // Пишем в кеш опкода
            op_cache <= i_data;
            pc <= pc + 1'b1;
            am <= 1'b0;
        
            // -----------------------
            /* ИНСТРУКЦИИ АЛУ */
            // -----------------------
            
            casex (opcode)
            
                // Indirect,X   (Непрямой,X)            ($FF,X)
                // -----------------------------------------------------
                8'bxxx_000_x1: t <= 4'h1;                
                
                // Zero Page    (Нуль-страница)         $FF
                // -----------------------------------------------------
                8'bxxx_001_xx, 
                8'b1xx_00x_00: t <= 4'h2;

                // Immediate    (Непосредственный)      #$FF
                // -----------------------------------------------------
                8'bxxx_010_x1: t <= 4'hC; // Перейти сразу к исполнению

                // Absolute     (Абсолютный 16)         $FFFF
                // -----------------------------------------------------
                8'bxxx_011_xx, 
                8'b001_000_00: t <= 4'h3;
                
                // Indirect,Y   (Непрямой),Y            ($FF),Y
                // -----------------------------------------------------
                8'bxxx_100_x1: 
                begin end
                
                // Zero Page,X  (Смещение 8 + X)        $FF,X
                // -----------------------------------------------------
                8'bxxx_101_xx: 
                begin end // + 4 ZPY
                
                // Absolute,Y   (Абсолютный 16 + Y)     $FFFF,Y
                // -----------------------------------------------------
                8'bxxx_110_x1, 
                8'b10x_111_1x: t <= 4'h4;

                // Absolute,X   (Абсолютный 16 + X)     $FFFF,X
                // -----------------------------------------------------
                8'bxxx_111_xx: t <= 4'h5;
                
                // Relative     (Условные переходы)     Метка (-128..127)
                // -----------------------------------------------------
                8'bxxx_100_00: 
                begin end
                
                // Implied      (Нет операндов)
                // -----------------------------------------------------
                default: 
                begin end

            endcase
        
        end
        
        /*
         * Чтение операндов
         */
        
        // Indirect,X
        4'h1: case (am)
            
            3'h0: begin am <= 3'h1; addr[15:0] <= {8'h00, i_data + x}; alt <= 1'b1; end // Перейти к этому адресу (Addr + X)
            3'h1: begin am <= 3'h2; tmp8 <= i_data; addr[7:0] <= addr[7:0] + 1'b1; end // Прочитать младший байт
            3'h2: begin t  <= 4'hC; addr <= {i_data, tmp8}; end // Проставить новый указатель для чтения операнда и переход к исполнению
        
        endcase

        // Zero Page
        4'h2: begin alt <= 1'b1; addr <= i_data; t <= 4'hC; end // Читать байт из указанной в ZP 
        
        // 3 - Absolute
        // 4 - Absolute,Y
        // 5 - Absolute,X
        4'h3, 4'h4, 4'h5: case (am)
        
            3'h0: begin am <= 3'h1; tmp8 <= i_data; pc <= pc + 1'b1; end // Читать младший байт
            3'h1: begin t  <= 4'hC; addr <= {i_data, tmp8} + (t == 4'h4 ? x : (t == 4'h5 ? y : 0)); pc <= pc + 1'b1; alt <= 1'b1; end // Старший байт [+X,Y]
        
        endcase

        /*
         * Исполнение опкодов
         */       
        
        4'hC: begin 
        
            // ---
        
        end

    endcase

end

endmodule
