`timescale 10ns / 1ns

module main;

// ---------------------------------------------------------------------

reg         clk;
always #0.5 clk         = ~clk;

initial begin clk = 1; #2000 $finish; end
initial begin $dumpfile("result.vcd"); $dumpvars(0, main); end

// ---------------------------------------------------------------------

endmodule
