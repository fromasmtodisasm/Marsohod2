/* 
 * Не находится в ведении копирайтов. Сделан, как кофе с утра.
 * Реклама: я кот, хозяин спит, лей вискаса, а то разодру обои.
 */
 
module z80(

    // О`клок
    input wire          clk,    /* 25 Мгц. Любой. */

    // Кот    #1 Порт
    output reg [15:0]   Ca,     /* Адрес памяти для считывания кода */
    input wire [7:0]    Ci,     /* Считанный код */
    
    // Данные #2 Порт
    output reg [15:0]   Da,     /* Для считывания данных */
    input wire [7:0]    Di,     /* Считанные данные */
    output reg [7:0]    Do,     /* Данные на запись */
    output reg          Dw      /* Сигнал записи */

);

// Методы адресации к Da
`define DA_PCI   3'b000
`define DA_BCDE  3'b001
`define DA_TINC  3'b010
`define DA_CIT   3'b011

// ---------------------------------------------------------------------
/* Основной набор регистров (8x8 = 256 бит) */
reg [7:0]  B; reg [7:0] C;
reg [7:0]  D; reg [7:0] E;
reg [7:0]  H; reg [7:0] L;
reg [7:0]  A; reg [7:0] F;
reg [15:0] IX;
reg [15:0] IY;
reg [15:0] SP;
reg [15:0] PC;
reg [ 7:0] I;   /* Прерывание */
reg [ 7:0] R;   /* Регенерация */
reg [ 1:0] IMODE;
reg        IFF1;
reg        IFF2;
reg        HALT;

/* Дополнительный набор. Регистры много занимают памяти в ПЛИС. */
reg [7:0] B_; reg [7:0] C_;
reg [7:0] D_; reg [7:0] E_;
reg [7:0] H_; reg [7:0] L_;
reg [7:0] A_; reg [7:0] F_;

/* Текущий регистр */
reg [2:0] Rq;   /* Запрос чтения */
reg [7:0] Rc;   /* Ответ чтения */

/* Для записи в регистр */
reg [2:0] Wn;   /* Номер регистра */
reg [7:0] Wo;   /* Значение */
reg       We;   /* Сигнал записи на следующем такте */

/* Префиксирование */
reg [1:0] Px;   /* Префиксировано 00 - HL; 01 - IX; 10 - IY; 11 - ?? */
reg [7:0] Hp;   /* Регистр H */
reg [7:0] Lp;   /* Регистр L */

// Состояние процессора
// ---------------------------------------------------------------------
reg [1:0] M_cycle;

// ---------------------------------------------------------------------

/* Инициализация регистров */
initial begin

    PC   = 16'h0000;
    SP   = 16'h0000;
    IX   = 16'h0000;
    IY   = 16'h0000;
    
    Rq   = 3'b000;
    Dw   = 1'b0;
    Px   = 2'b00;
    T    = 8'h00;
    
    /* Специальные регистры */
    IMODE = 2'b00;
    IFF1  = 1'b0;
    IFF2  = 1'b0;
    HALT  = 1'b0;
    {I, R} = {8'h00, 8'h00};
    
    M_cycle = 1'b0;
    
    //                                      B      C      D      E      H      L      A      F
    {B,  C,  D,  E,  H,  L,  A,  F } = {8'h02, 8'h00, 8'h01, 8'h05, 8'h05, 8'h12, 8'h41, 8'h00};
    {B_, C_, D_, E_, H_, L_, A_, F_} = {8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFA, 8'h00};

end

// Эмуляция микрокода
// ---------------------------------------------------------------------

reg [1:0]   mPCinc;           /* Увеличить PC + mPCinc на следующем такте */

reg         mPCrel;           /* Если =1, переход на jmpRel */
reg         mPCjmp;           /* Признак, что есть переход на PCtmp */
reg [15:0]  PCrel;            /* Вычисление относительн PC перехода 8 бит */

reg         iMC;              /* Увеличить M_cycle */
reg         mEXAF;            /* На следующем такте развернуть AF, AF' */
reg         mBDec;            /* B = B - 1 */

reg [1:0]   We16;             /* Запись в 16-битный регистр Wn[1:0] */
reg [1:0]   mT;               /* Действия с регистром T */
reg [15:0]  T;                /* Временное значение */
reg [2:0]   DaS;              /* Источник Da */

reg [15:0]  refDEBC;

/* Кеш опкода между M_cycle */
reg [7:0]   opcache;      

/* Источник опкода */
wire [7:0]  opcode = (M_cycle == 1'b0) ? Ci : opcache;  

/* Проверка условий */
wire [3:0]  condition = { F[7], F[2], F[6], F[0] };

/* Для двухбайтовой записи в память или из памяти */
wire [15:0] Tinc = T + 1'b1;

/* Частично считанные данные */
wire [15:0] DiT  = {Di[7:0], T[7:0]};

// ---------------------------------------------------------------------

always @* begin

    Ca          = PC;
    DaS         = `DA_PCI;
    Dw          = 1'b0;
    DaS         = 1'b0;
    
    /* Секция переходов */
    iMC         = 1'b0;
    mPCinc      = 2'b01;
    mPCjmp      = 1'b0;
    mPCrel      = 1'b0;      
     PCrel      = PC + {{8{Di[7]}}, Di[7:0]} + 2'h2;
        
    /* Запись в регистры */
    mEXAF       = 1'b0;
    mBDec       = 1'b0;
    We16        = 2'b00;
    mT          = 2'b00;
    We          = 1'b0;
    Wn          = opcode[5:3];

    casex (opcode)
            
        // 1T EX AF, AF'
        8'b00_001_000: mEXAF = 1'b1; 
        
        // 1T DJNZ *
        8'b00_010_000: {mBDec, mPCinc, mPCrel} = {1'b1, 2'b10, (B != 8'h00) };

        // 1T JR *
        8'b00_011_000: {mPCrel} = {1'b1};
        
        // 1T JR {NC, C, NZ, Z}, *
        8'b00_1xx_000: {mPCinc, mPCrel} = {2'b10, condition[ opcode[4] ] == opcode[3] };
        
        // 2T LD r16, **
        8'b00_xx0_001: case (M_cycle)
        
            /* Запись из Di -> T[7:0], PC += 2 */
            1'b0: {iMC, mT} = {1'b1, 2'b01};
            
            /* Запись {Di, T[7:0]} -> r16 */
            1'b1: {We16, Wn[1:0]} = {2'b01, opcode[5:4]};
        
        endcase
        
        // -------------------------------------------------------------
        
        
        // ADD HL, r16
        // 8'b00_xx1_001:  ----------
        
        // 2T LD (r16), A :: Запись в память (BC|DE)
        8'b00_0x0_010: case (M_cycle)
        
            /* Подготовка шины к записи */
            1'b0: {iMC, mPCinc} <= {1'b1, 2'b01};
        
            /* Запись на шину Da */
            1'b1: {DaS, mPCinc, Dw, Do} <= {3'b001, 2'b00, 1'b1, A};

        endcase
        
        // 2T LD A, (r16) :: Чтение из памяти (BC|DE)
        8'b00_0x1_010: case (M_cycle)
        
            /* Ожидание появления валидных данных на шине Da */
            1'b0: {iMC, mPCinc} <= {1'b1, 2'b00};

            /* Запись данных в регистр с шины Da */
            1'b1: {DaS, We, Wn, Wo} <= {3'b001, 1'b1, 3'b111, Di};
            
        endcase
        
        // 4T LD (**), HL
        8'b00_100_010: case (M_cycle)
        
            /* Записать Di -> T[7:0], PC += 2 */
            1'b0: {iMC, mT, mPCinc} = {1'b1, 2'b01, 2'b10};

            /* Установка адреса и запись L. Запись Ci -> T[15:8] */
            1'b1: {iMC, mT, DaS, mPCinc} = {1'b1, 2'b10, 3'b011, 2'b00};
            
            /* Запись HL в память */
            2'h2: {iMC, DaS, Dw, Do, mPCinc} = {1'b1, 3'b011, 1'b1, L, 2'b00};
            2'h3: {DaS, Dw, Do} = {3'b010, 1'b1, H};
        
        
        // LD HL, (**)
        8'b00_101_010: case (M_cycle)
        
            /* Записать Di -> T[7:0], PC += 2 */
            1'b0: {iMC, mT, mPCinc}     = {1'b1, 2'b01, 2'b10};
            1'b1: {iMC, mT, DaS, mPCinc} = {1'b1, 2'b10, 3'b011, 2'b00 };
            //2'h2: {Ca, Da, nWe16, Wn[1:0]} = {Tinc, T, 2'b10, 2'b10};
        
        endcase
        
        endcase
    
    endcase

    /* Источник Da */
    case (DaS)
    
        `DA_BCDE: Da = opcode[4] ? {D,E} : {B,C};
        `DA_TINC: Da = T + 1'b1;
        `DA_CIT:  Da = {Ci[7:0], T[7:0]};
        default:  Da = PC + 1'b1;
    
    endcase
    
end


// Тактирование. Основная логика
// ---------------------------------------------------------------------

always @(posedge clk) begin

    /* Переходы */
    PC <= mPCrel ? PCrel :  PC + mPCinc;
    
    /* Обработка T16 */
    case (mT)
    
        2'b01: T[7:0]  <= Di;
        2'b10: T[15:8] <= Ci;
        
    endcase    
        
    /* Запись опкода в кеш */
    if (M_cycle == 1'b0)
        opcache <= Ci;

    /* Есть следующий опкод */
    if (iMC) begin
        
        M_cycle <= M_cycle + 1'b1;
        
    end else begin /* Финализация. Регистр регенерации. */
    
        M_cycle <= 1'b0;
        R[6:0]  <= R[6:0] + 1'b1;
        
    end
    
end


/* Чтение из регистров */
// ---------------------------------------------------------------------

always @(Rq, Px, mEXAF) begin

    case (Px)
        2'b00: begin Hp = H;        Lp = L; end
        2'b01: begin Hp = IX[15:8]; Lp = IX[7:0]; end
        2'b10: begin Hp = IY[15:8]; Lp = IY[7:0]; end
    endcase
        
    /* Другие инструкции */
    case (Rq)
        
        3'b000: Rc = B;  3'b001: Rc = C;
        3'b010: Rc = D;  3'b011: Rc = E;
        3'b100: Rc = Hp; 3'b101: Rc = Lp;
        3'b110: Rc = Di; 3'b111: Rc = A; 
    
    endcase

end

/* Запись в регистры */
// ---------------------------------------------------------------------

always @(posedge clk) begin

    /* Команда EX AF, AF' */
    if (mEXAF) {A, A_, F, F_} <= {A_, A, F_, F};
    
    /* Уменьшение B = B - 1 */
    else if (mBDec) B <= B - 1'b1;    
    
    /* Запись в регистр 16 бит из памяти {Di, T[7:0]} */
    else if (We16 == 2'b01) begin
    
        case (Wn[1:0])
        
            2'b00: {B, C} <= DiT;
            2'b01: {D, E} <= DiT;
            2'b10: {H, L} <= DiT;
            2'b11: SP     <= DiT;

        endcase
    
    end
        
    /* Регистр */
    else if (We) begin

        case (Wn)
            3'b000: B <= Wo;  3'b001: C <= Wo;
            3'b010: D <= Wo;  3'b011: E <= Wo;
            3'b100: case (Px) 2'b00:  H <= Wo; 2'b01: IX[15:8] <= Wo; 2'b10: IY[15:8] <= Wo; endcase
            3'b101: case (Px) 2'b00:  L <= Wo; 2'b01: IX[ 7:0] <= Wo; 2'b10: IY[ 7:0] <= Wo; endcase
            // 3'b110: /* Запись в память обрабатывается отдельно */ begin Dw <= We; Do <= Wo;  end
            3'b111: A <= Wo;
        endcase

    end
    
    /* Флаги */
    // ... 
    
    // Другое (SP и прочее)

end

endmodule
