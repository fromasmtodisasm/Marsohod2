/* 
 * Не находится в ведении копирайтов. Сделан, как кофе с утра.
 * Реклама: я кот, хозяин спит, лей вискаса, а то разодру обои.
 */
 
module z80(

    // О`клок
    input wire          clk,    /* 25 Мгц. Любой. */

    // Кот    #1 Порт
    output reg [15:0]   PC,     /* Адрес памяти для считывания кода */
    input wire [7:0]    Ci,     /* Считанный код */
    
    // Данные #2 Порт
    output reg [15:0]   Da,     /* Для считывания данных */
    input wire [7:0]    Di,     /* Считанные данные */
    output reg [7:0]    Do,     /* Данные на запись */
    output reg          Dw      /* Сигнал записи */

);

// ---------------------------------------------------------------------
/* Основной набор регистров (8x8 = 256 бит) */
reg [7:0]  B; reg [7:0] C;
reg [7:0]  D; reg [7:0] E;
reg [7:0]  H; reg [7:0] L;
reg [7:0]  A; reg [7:0] F;
reg [15:0] IX;
reg [15:0] IY;
reg [15:0] SP;

/* Дополнительный набор. Регистры много занимают памяти в ПЛИС. */
reg [7:0] B_; reg [7:0] C_;
reg [7:0] D_; reg [7:0] E_;
reg [7:0] H_; reg [7:0] L_;
reg [7:0] A_; reg [7:0] F_;

/* Если = 0, то указывает на набор 0, иначе на 1 */
reg       Bank;

/* Текущий регистр */
reg [2:0] Rq;   /* Запрос */
reg [7:0] Rc;   /* Ответ  */
reg [1:0] Px;   /* Префиксировано 00 - HL; 01 - IX; 10 - IY; 11 - ?? */
reg [7:0] Hp;   /* Регистр H (префикс может) */
reg [7:0] Lp;   /* Регистр L (префикс может) */

// ---------------------------------------------------------------------

/* Инициализация регистров */
initial begin

    PC   = 16'h0000;
    SP   = 16'h0000;
    IX   = 16'h0000;
    IY   = 16'h0000;
    
    Rq   = 3'b000;
    Px   = 2'b00;
    Bank = 1'b0;
    
    {B,  C,  D,  E,  H,  L,  A,  F} = 64'h0;
    {B_, C_, D_, E_, H_, L_, A_, F_} = 64'h0;

end

// Тактирование. Основная логика.
// ---------------------------------------------------------------------

always @(posedge clk) begin

    PC <= PC + 1'b1;

end

// Выборка регистра
// ---------------------------------------------------------------------

always @(Px, Bank, Rq) begin

    case (Px)
        2'b00: begin Hp = Bank ? H_ : H;
                     Lp = Bank ? L_ : L; end
        2'b01: begin Hp = IX[15:8]; Lp = IX[7:0]; end
        2'b10: begin Hp = IY[15:8]; Lp = IY[7:0]; end
    endcase

    case ({Bank, Rq})
        
        /* Банк 0 */
        4'b0_000: Rc = B;  4'b0_001: Rc = C;
        4'b0_010: Rc = D;  4'b0_011: Rc = E;
        4'b0_100: Rc = Hp; 4'b0_101: Rc = Lp;
        4'b0_110: Rc = Di; /* (HL,IX,IY) */
        4'b0_111: Rc = A; 
    
        /* Банк 1 */
        4'b1_000: Rc = B_; 4'b1_001: Rc = C_;
        4'b1_010: Rc = D_; 4'b1_011: Rc = E_;
        4'b1_100: Rc = Hp; 4'b1_101: Rc = Lp;
        4'b1_110: Rc = Di; /* (HL,IX,IY) */
        4'b1_111: Rc = A_;

    endcase

end

endmodule
